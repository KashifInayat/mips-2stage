module main(
input clk,
input rst,
input interrupt1,
input [7:0]  key_code1,
output  [31:0]for_display,
output  [31:0]for_display1,
output [9:0] count_out

);
//controller
wire jal;
wire lui;
wire lli;
wire ctl1;
wire ctl2;
wire ctl3;
wire ctl4;
wire ctl5;
wire ctl7;
wire ctl8;
wire ctl9;
//counter
//wire [9:0] count_out;//counter output
//pm
wire p_enbl_a;
wire p_enbl_b;
wire  [31:0] inst_a;
wire [31:0] inst_b;
reg [31:0] inst_out;//pm output
//reg file
reg [31:0] dm_alu_out;
reg [15:0] lsb_reg_in;
reg [15:0] msb_reg_in;
wire [31:0] bt0;
wire [31:0]reg_out1;//reg out 1
wire [31:0]reg_out2;//reg out 2
/////////Memory Map register////////
reg [31:0] r_map;
wire map_e;
reg map_and;
reg [31:0] dm_out;
//dm nd mux
wire d_enbl_a;
wire d_enbl_b;
wire  [31:0] dm_a;
wire [31:0] dm_b;
reg [9:0]addr_in;
reg [31:0] dm_out1;//dm output
//alu
reg [31:0] data2_alu_in;
wire [31:0] data_alu_out;
//Pipelining Register's and Mux's.
reg [31:0]inst_r_1;
reg [31:0]reg_d01;
reg ctl2_1;
reg ctl7_1;
reg ctl1_1;
reg lui_1;
reg lli_1;
reg [31:0]mux_d02;
reg [31:0]inst_r_2;
reg [31:0]mux_alu_o;
reg ctl7_2;
reg ctl1_2;
reg lui_2;
reg lli_2;
//forwarding Muxes nd Select lines(read after write)
reg [31:0] fw_d1;
wire sel_md1; 
reg [31:0] fw_d2;
wire sel_md2;
//forwarding Mux nd Select line(write after write)
wire sel_dm;
reg [31:0] fw_dm;
//Controller
control_unit inst(
.clk(clk),
.rst(rst),
.bt0(bt0),
.opcode(inst_out[31:27]),
.jal(jal),
.lui(lui),
.lli(lli),
.ctl1(ctl1),
.ctl2(ctl2),
.ctl3(ctl3),
.ctl4(ctl4),
.ctl5(ctl5),
.ctl7(ctl7),
.ctl8(ctl8),
.ctl9(ctl9)
);
//counter
pc inst1(
.clk(clk),
.rst(rst),
.sel_m1(ctl4),
.sel_m2(ctl5),
.inst_pm(inst_out[9:0]),
.reg_out(reg_out1[9:0]),
.count(count_out)
);

//Program Memory 
assign p_enbl_a = (count_out[9:8]==2'b00);
assign p_enbl_b = (count_out[9:8]==2'b01);
//  RAMB16_S36 : In order to incorporate this function into the design,
//   Verilog   : the following instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB16_S36_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB16_S36: 512 x 32 + 4 Parity bits Single-Port RAM
   //             Spartan-3E
   // Xilinx HDL Language Template, version 12.1

RAMB16_S36 #(
      .INIT(36'h000000000),  // Value of output RAM registers at startup
      .SRVAL(36'h000000000), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 127
      .INIT_00(256'h21c00005_21c00004_21c00003_21c00002_21c00001_21c00000_f0000000_4800024a),
      .INIT_01(256'h21c0000d_21c0000c_21c0000b_21c0000a_21c00009_21c00008_21c00007_21c00006),
      .INIT_02(256'h480003e8_21c00014_21c00013_21c00012_21c00011_21c00010_21c0000f_21c0000e),
      .INIT_03(256'h21c0001b_21c0001a_21c00019_21c00018_21c00017_21c00016_21c00015_f0000000),
      .INIT_04(256'h21c00023_21c00022_21c00021_21c00020_21c0001f_21c0001e_21c0001d_21c0001c),
      .INIT_05(256'hf0000000_480003d1_21c00029_21c00028_21c00027_21c00026_21c00025_21c00024),
      .INIT_06(256'h21c00031_21c00030_21c0002f_21c0002e_21c0002d_21c0002c_21c0002b_21c0002a),
      .INIT_07(256'h21c00039_21c00038_21c00037_21c00036_21c00035_21c00034_21c00033_21c00032),
      .INIT_08(256'h21c0003f_f0000000_480003ba_21c0003e_21c0003d_21c0003c_21c0003b_21c0003a),
      .INIT_09(256'h21c00047_21c00046_21c00045_21c00044_21c00043_21c00042_21c00041_21c00040),
      .INIT_0A(256'h21c0004f_21c0004e_21c0004d_21c0004c_21c0004b_21c0004a_21c00049_21c00048),
      .INIT_0B(256'h21c00056_21c00054_f0000000_480003a3_21c00053_21c00052_21c00051_21c00050),
      .INIT_0C(256'h21c0005e_21c0005d_21c0005c_21c0005b_21c0005a_21c00059_21c00058_21c00057),
      .INIT_0D(256'h21c00066_21c00065_21c00064_21c00063_21c00062_21c00061_21c00060_21c0005f),
      .INIT_0E(256'h21c0006c_21c0006b_21c0006a_21c00069_f0000000_4800038d_21c00068_21c00067),
      .INIT_0F(256'h21c00074_21c00073_21c00072_21c00071_21c00070_21c0006f_21c0006e_21c0006d),
      // Address 128 to 255
      .INIT_10(256'h21c0007c_21c0007b_21c0007a_21c00079_21c00078_21c00077_21c00076_21c00075),
      .INIT_11(256'h21c00082_21c00081_21c00080_21c0007f_21c0007e_f0000000_48000376_21c0007d),
      .INIT_12(256'h21c0008a_21c00089_21c00088_21c00087_21c00086_21c00085_21c00084_21c00083),
      .INIT_13(256'h21c00092_21c00091_21c00090_21c0008f_21c0008e_21c0008d_21c0008c_21c0008b),
      .INIT_14(256'h21c00098_21c00097_21c00096_21c00095_21c00094_21c00093_f0000000_4800035f),
      .INIT_15(256'h21c000a0_21c0009f_21c0009e_21c0009d_21c0009c_21c0009b_21c0009a_21c00099),
      .INIT_16(256'h48000348_21c000a7_21c000a6_21c000a5_21c000a4_21c000a3_21c000a2_21c000a1),
      .INIT_17(256'h21c000ae_21c000ad_21c000ac_21c000ab_21c000aa_21c000a9_21c000a8_f0000000),
      .INIT_18(256'h21c000b6_21c000b5_21c000b4_21c000b3_21c000b2_21c000b1_21c000b0_21c000af),
      .INIT_19(256'hf0000000_48000331_21c000bc_21c000bb_21c000ba_21c000b9_21c000b8_21c000b7),
      .INIT_1A(256'h21c000c4_21c000c3_21c000c2_21c000c1_21c000c0_21c000bf_21c000be_21c000bd),
      .INIT_1B(256'h21c000cc_21c000cb_21c000ca_21c000c9_21c000c8_21c000c7_21c000c6_21c000c5),
      .INIT_1C(256'h21c000d4_21c000d3_21c000d2_21c000d1_21c000d0_21c000cf_21c000ce_21c000cd),
      .INIT_1D(256'h21c000dc_21c000db_21c000da_21c000d9_21c000d8_21c000d7_21c000d6_21c000d5),
      .INIT_1E(256'h21c000e4_21c000e3_21c000e2_21c000e1_21c000e0_21c000df_21c000de_21c000dd),
      .INIT_1F(256'h21c000ea_21c000e9_21c000e8_21c000e7_21c000e6_21c000e5_f0000000_48000307),
      // Address 256 to 383
      .INIT_20(256'h21c000f2_21c000f1_21c000f0_21c000ef_21c000ee_21c000ed_21c000ec_21c000eb),
      .INIT_21(256'h21c000fa_21c000f9_21c000f8_21c000f7_21c000f6_21c000f5_21c000f4_21c000f3),
      .INIT_22(256'h21c00102_21c00101_21c00100_21c000ff_21c000fe_21c000fd_21c000fc_21c000fb),
      .INIT_23(256'h21c0010a_21c00109_21c00108_21c00107_21c00106_21c00105_21c00104_21c00103),
      .INIT_24(256'h21c00110_21c0010f_21c0010e_21c0010d_f0000000_480002dd_21c0010c_21c0010b),
      .INIT_25(256'h21c00118_21c00117_21c00116_21c00115_21c00114_21c00113_21c00112_21c00111),
      .INIT_26(256'h21c00120_21c0011f_21c0011e_21c0011d_21c0011c_21c0011b_21c0011a_21c00119),
      .INIT_27(256'h21c00128_21c00127_21c00126_21c00125_21c00124_21c00123_21c00122_21c00121),
      .INIT_28(256'h21c00130_21c0012f_21c0012e_21c0012d_21c0012c_21c0012b_21c0012a_21c00129),
      .INIT_29(256'h21c00136_21c00135_f0000000_480002b3_21c00134_21c00133_21c00132_21c00131),
      .INIT_2A(256'h21c0013e_21c0013d_21c0013c_21c0013b_21c0013a_21c00139_21c00138_21c00137),
      .INIT_2B(256'h21c00146_21c00145_21c00144_21c00143_21c00142_21c00141_21c00140_21c0013f),
      .INIT_2C(256'h21c0014e_21c0014d_21c0014c_21c0014b_21c0014a_21c00149_21c00148_21c00147),
      .INIT_2D(256'h21c00156_21c00155_21c00154_21c00153_21c00152_21c00151_21c00150_21c0014f),
      .INIT_2E(256'hf0000000_48000289_21c0015c_21c0015b_21c0015a_21c00159_21c00158_21c00157),
      .INIT_2F(256'h21c00164_21c00163_21c00162_21c00161_21c00160_21c0015f_21c0015e_21c0015d),
      // Address 384 to 511
      .INIT_30(256'h21c0016c_21c0016b_21c0016a_21c00169_21c00168_21c00167_21c00166_21c00165),
      .INIT_31(256'h21c00174_21c00173_21c00172_21c00171_21c00170_21c0016f_21c0016e_21c0016d),
      .INIT_32(256'h21c0017c_21c0017b_21c0017a_21c00179_21c00178_21c00177_21c00176_21c00175),
      .INIT_33(256'h21c00184_21c00183_21c00182_21c00181_21c00180_21c0017f_21c0017e_21c0017d),
      .INIT_34(256'h21c0018a_21c00189_21c00188_21c00187_21c00186_21c00185_f0000000_4800025f),
      .INIT_35(256'h21c00192_21c00191_21c00190_21c0018f_21c0018e_21c0018d_21c0018c_21c0018b),
      .INIT_36(256'h21c0019a_21c00199_21c00198_21c00197_21c00196_21c00195_21c00194_21c00193),
      .INIT_37(256'h21c001a2_21c001a1_21c001a0_21c0019f_21c0019e_21c0019d_21c0019c_21c0019b),
      .INIT_38(256'h21c001aa_21c001a9_21c001a8_21c001a7_21c001a6_21c001a5_21c001a4_21c001a3),
      .INIT_39(256'h21c001b0_21c001af_21c001ae_21c001ad_f0000000_48000235_21c001ac_21c001ab),
      .INIT_3A(256'h21c001b8_21c001b7_21c001b6_21c001b5_21c001b4_21c001b3_21c001b2_21c001b1),
      .INIT_3B(256'h21c001c0_21c001bf_21c001be_21c001bd_21c001bc_21c001bb_21c001ba_21c001b9),
      .INIT_3C(256'h21c001c8_21c001c7_21c001c6_21c001c5_21c001c4_21c001c3_21c001c2_21c001c1),
      .INIT_3D(256'h21c001d0_21c001cf_21c001ce_210001cd_21c001cc_21c001cb_21c001ca_21c001c9),
      .INIT_3E(256'h21c001d6_21c001d5_f0000000_4800020b_21c001d4_21c001d3_21c001d2_21c001d1),
      .INIT_3F(256'h21c001de_210001dd_21c001dc_21c001db_21c001da_21c001d9_21c001d8_21c001d7),

      // The next set of INITP_xx are for the parity bits
      // Address 0 to 127
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 128 to 255
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 256 to 383
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 384 to 511
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) PM_inst1 (
      .DO(inst_a),      // 32-bit Data Output
      .DOP(),    // 4-bit parity Output
      .ADDR(count_out[8:0]),  // 9-bit Address Input
      .CLK(clk),    // Clock
      .DI(32'd0),      // 32-bit Data Input
      .DIP(4'd0),    // 4-bit parity Input
      .EN(p_enbl_a),      // RAM Enable Input
      .SSR(rst),    // Synchronous Set/Reset Input
      .WE(1'd0)       // Write Enable Input
   );

// End of RAMB16_S36_inst instantiation
//Program Memory 

//  RAMB16_S36 : In order to incorporate this function into the design,
//   Verilog   : the following instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB16_S36_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB16_S36: 512 x 32 + 4 Parity bits Single-Port RAM
   //             Spartan-3E
   // Xilinx HDL Language Template, version 12.1

RAMB16_S36 #(
      .INIT(36'h000000000),  // Value of output RAM registers at startup
      .SRVAL(36'h000000000), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 127
      .INIT_00(256'h21c001e6_21c001e5_21c001e4_21c001e3_21c001e2_21c001e1_21c001e0_21c001df),
      .INIT_01(256'h21c001ee_210001ed_21c001ec_21c001eb_21c001ea_21c001e9_21c001e8_21c001e7),
      .INIT_02(256'h21c001f6_21c001f5_21c001f4_21c001f3_21c001f2_21c001f1_21c001f0_21c001ef),
      .INIT_03(256'hf0000000_480002e1_21c001fc_21c001fb_21c001fa_21c001f9_21c001f8_21c001f7),
      .INIT_04(256'h21c00204_21c00203_21c00202_21c00201_21c00200_210001ff_21c001fe_210001fd),
      .INIT_05(256'h21c0020c_21c0020b_21c0020a_21c00209_21c00208_21c00207_21c00206_21c00205),
      .INIT_06(256'h21c00214_21c00213_21c00212_21c00211_21c00210_2100020f_21c0020e_2100020d),
      .INIT_07(256'h21c0021c_21c0021b_21c0021a_21c00219_21c00218_21c00217_21c00216_21c00215),
      .INIT_08(256'h21c00224_21c00223_21c00222_21c00221_21c00220_2100021f_21c0021e_2100021d),
      .INIT_09(256'h00000000_00000000_00000000_480003fe_224002bc_00000000_f0000000_480001b7),
      .INIT_0A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 128 to 255
      .INIT_10(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_11(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_12(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_13(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_14(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_15(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_16(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_17(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_18(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_19(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 256 to 383
      .INIT_20(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_21(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_22(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_23(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_24(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_25(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_26(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_27(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_28(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_29(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 384 to 511
      .INIT_30(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_31(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_32(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_33(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_34(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_35(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_36(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_37(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_38(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_39(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),

      // The next set of INITP_xx are for the parity bits
      // Address 0 to 127
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 128 to 255
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 256 to 383
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 384 to 511
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) 
   PM_inst2 (
      .DO(inst_b),      // 32-bit Data Output
      .DOP(),    // 4-bit parity Output
      .ADDR(count_out[8:0]),  // 9-bit Address Input
      .CLK(clk),    // Clock
      .DI(32'd0),      // 32-bit Data Input
      .DIP(4'd0),    // 4-bit parity Input
      .EN(p_enbl_b),      // RAM Enable Input
      .SSR(rst),    // Synchronous Set/Reset Input
      .WE(1'd0)       // Write Enable Input
   );

// End of RAMB16_S36_inst instantiation
    always@(*)
  begin
  case(p_enbl_b)
    1'd0: inst_out=inst_a;
    1'd1: inst_out=inst_b;
    
  endcase
end
///////////End Of Pm
//MUXES for reg 
    always@(*)
  begin
  case(ctl2_1)
    1'd0: dm_alu_out=data_alu_out;
    1'd1: dm_alu_out=dm_out;
    
  endcase
end

//Pipelining before Reg File Written Side

//2nd Inst register 
always@(posedge clk)
   begin
     if(rst)
      inst_r_2 <=#1 0;
     else
       inst_r_2 <=#1 inst_r_1;
   end

//Reg File MUX of (ALU Out +DM Out)+ Instruction data Register(written Side)
always@(posedge clk)
   begin
     if(rst)
      mux_alu_o <= #1 0;//register
     else
       mux_alu_o <= #1 dm_alu_out;//register
   end   

// 2nd Register For CTL7
always@(posedge clk)
   begin
     if(rst)
      ctl7_2 <= #1 0;
     else
      ctl7_2 <= #1 ctl7_1;
   end  

// 2nd Register For CTL1
always@(posedge clk)
   begin
     if(rst)
      ctl1_2 <= #1 0;
     else
      ctl1_2 <= #1 ctl1_1;
   end 
   
// 2nd Register For lui
always@(posedge clk)
   begin
     if(rst)
      lui_2 <= #1 0;
     else
      lui_2 <= #1 lui_1;
   end 
   
// 2nd Register For lli
always@(posedge clk)
   begin
     if(rst)
      lli_2 <= #1 0;
     else
      lli_2 <= #1 lli_1;
   end 
// end of Pipelining before Reg File Written Side

  //for 16 lsb reg in
  always@(*)
  begin
  case(ctl7_2)
    1'd0: lsb_reg_in=mux_alu_o[15:0];
    1'd1: lsb_reg_in=inst_r_2[15:0];
    
  endcase
end
//for 16 msb reg in
  always@(*)
  begin
  case(ctl7_2)
    1'd0: msb_reg_in=mux_alu_o[31:16];
    1'd1: msb_reg_in=inst_r_2[15:0];
    
  endcase
end		
//reg File
reg_file inst2(
  .clk(clk),
	.rd_addr1(inst_out[21:17]),
	.rd_addr2(inst_out[16:12]),
	.wr_addr(inst_r_2[26:22]),
	.wr_data1(lsb_reg_in),
  .wr_data2(msb_reg_in),
	.count_out(count_out),
	.jal(jal),
	.wr_en(ctl1_2),
	.wr_en_upr(lui_2),
	.wr_en_lwr(lli_2),
	.rd_data1(reg_out1),
	.rd_data2(reg_out2),
	.for_display1(for_display1),
	.for_display(for_display),
	.bt(bt0)
		);
//MUX for dm
  always@(*)
  begin
  case(ctl9)
    1'd0: addr_in=inst_out[9:0];
    1'd1: addr_in=reg_out2[9:0];
    
  endcase
end				
//Mux for forwarding (write after write)				
//Mux dm_data_ Select Line
assign sel_dm=(inst_out[21:17]==inst_r_2[26:22]);
//Mux dm_data  
  always@(*)
  begin
  case(sel_dm)
    1'd0: fw_dm=reg_out1;
    1'd1: fw_dm=mux_alu_o;
    
  endcase
end
////////////////////dm///////////////

assign d_enbl_a = (addr_in[9:8]==2'b00);
assign d_enbl_b = (addr_in[9:8]==2'b01);
//  RAMB16_S36 : In order to incorporate this function into the design,
//   Verilog   : the following instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB16_S36_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

// RAMB16_S36: 512 x 32 + 4 Parity bits Single-Port RAM
//             Spartan-3E
// Xilinx HDL Language Template, version 12.1
RAMB16_S36 #(
      .INIT(36'h000000000),  // Value of output RAM registers at startup
      .SRVAL(36'h000000000), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 127
      .INIT_00(256'h0000023E_0000023A_000001EF_000001E9_000001A0_00000198_00000151_00000147),
      .INIT_01(256'h000003C9_0000037E_0000037A_0000032D_0000032B_000002DC_0000028D_0000028B),
      .INIT_02(256'h000001B1_0000016A_00000160_00000471_00000467_00000420_00000418_000003CF),
      .INIT_03(256'h000002F5_000002A6_000002A4_00000257_00000253_00000208_00000202_000001B9),
      .INIT_04(256'h00000439_00000431_000003E8_000003E2_00000397_00000393_00000346_00000344),
      .INIT_05(256'h00000221_0000021B_000001D2_000001CA_00000183_00000179_0000048A_00000480),
      .INIT_06(256'h000003AC_0000035F_0000035D_0000030E_000002BF_000002BD_00000270_0000026C),
      .INIT_07(256'h00000737_000004A2_00000499_00000452_0000044A_00000401_000003FB_000003B0),
      .INIT_08(256'h0000087B_0000082E_0000082A_000007DF_000007D9_00000790_00000788_00000741),
      .INIT_09(256'h000009BF_000009B9_0000096E_0000096A_0000091D_0000091B_000008CC_0000087D),
      .INIT_0A(256'h000007A9_000007A1_0000075A_00000750_00000A60_00000A57_00000A10_00000A08),
      .INIT_0B(256'h00000934_000008E5_00000896_00000894_00000847_00000843_000007F8_000007F2),
      .INIT_0C(256'h00000A70_00000A29_00000A21_000009D8_000009D2_00000987_00000983_00000936),
      .INIT_0D(256'h0000085C_00000811_0000080B_000007C2_000007BA_00000773_00000769_00000A79),
      .INIT_0E(256'h000009A0_0000099C_0000094F_0000094D_000008FE_000008AF_000008AD_00000860),
      .INIT_0F(256'h00000D31_00000D27_00000A92_00000A89_00000A42_00000A3A_000009F1_000009EB),
      // Address 128 to 255
      .INIT_10(256'h00000E6D_00000E6B_00000E1E_00000E1A_00000DCF_00000DC9_00000D80_00000D78),
      .INIT_11(256'h00000FF8_00000FAF_00000FA9_00000F5E_00000F5A_00000F0D_00000F08_00000EBC),
      .INIT_12(256'h00000DE2_00000D99_00000D91_00000D4A_00000D40_00001050_00001047_00001000),
      .INIT_13(256'h00000F26_00000F24_00000ED5_00000E86_00000E84_00000E37_00000E33_00000DE8),
      .INIT_14(256'h00001069_00001060_0001019_000001011_00000FC8_00000FC2_00000F77_00000F73),
      .INIT_15(256'h00000E50_00000E4C_00000E01_00000DFB_00000DB2_00000DAA_00000D63_00000D59),
      .INIT_16(256'h00000FDB_00000F90_00000F8C_00000F3F_00000F3D_00000EEE_00000E9F_00000E9D),
      .INIT_17(256'h00000149_00000148_00000147_00001082_00001079_00001032_0000102A_00000FE1),
      .INIT_18(256'h00000151_00000150_0000014F_0000014E_0000014D_0000014C_0000014B_0000014A),
      .INIT_19(256'h00000291_00000287_00000241_00000237_000001F1_000001E7_000001A1_00000197),
      .INIT_1A(256'h000003D1_000003C7_00000381_00000377_00000331_00000327_000002E1_000002D7),
      .INIT_1B(256'h0000046C_0000046B_0000046A_00000469_00000468_00000467_00000421_00000417),
      .INIT_1C(256'h00000162_00000161_00000160_00000471_00000470_0000046F_0000046E_0000046D),
      .INIT_1D(256'h0000016A_00000169_00000168_00000167_00000166_00000165_00000164_00000163),
      .INIT_1E(256'h000002AA_000002A0_0000025A_00000250_0000020A_00000200_000001BA_000001B0),
      .INIT_1F(256'h000003EA_000003E0_0000039A_00000390_0000034A_00000340_000002FA_000002F0),
      // Address 256 to 383
      .INIT_20(256'h00000485_00000484_00000483_00000482_00000481_00000480_0000043A_00000430),
      .INIT_21(256'h0000017B_0000017A_00000179_0000048A_00000489_00000488_00000487_00000486),
      .INIT_22(256'h00000183_00000182_00000181_00000180_0000017F_0000017E_0000017D_0000017C),
      .INIT_23(256'h000002C3_000002B9_00000273_00000269_00000223_00000219_000001D3_000001C9),
      .INIT_24(256'h00000403_000003F9_000003B3_000003A9_00000363_00000359_00000313_00000309),
      .INIT_25(256'h0000049E_0000049D_0000049C_0000049B_0000049A_00000499_00000453_00000449),
      .INIT_26(256'h00000739_00000738_00000737_000004A3_000004A2_000004A1_000004A0_0000049F),
      .INIT_27(256'h00000741_00000740_0000073F_0000073E_0000073D_0000073C_0000073B_0000073A),
      .INIT_28(256'h00000881_00000877_00000831_00000827_000007E1_000007D7_00000791_00000787),
      .INIT_29(256'h000009C1_000009B7_00000971_00000967_00000921_00000917_000008D1_000008C7),
      .INIT_2A(256'h00000A5C_00000A5B_00000A5A_00000A59_00000A58_00000A57_00000A11_00000A07),
      .INIT_2B(256'h00000752_00000751_00000750_00000A61_00000A60_00000A5F_00000A5E_00000A5D),
      .INIT_2C(256'h0000075A_00000759_00000758_00000757_00000756_00000755_00000754_00000753),
      .INIT_2D(256'h0000089A_00000890_0000084A_00000840_000007FA_000007F0_000007AA_000007A0),
      .INIT_2E(256'h000009DA_000009D0_0000098A_00000980_0000093A_00000930_000008EA_000008E0),
      .INIT_2F(256'h00000A75_00000A74_00000A73_00000A72_00000A71_00000A70_00000A2A_00000A20),
      // Address 384 to 511
      .INIT_30(256'h0000076B_0000076A_00000769_00000A7A_00000A79_00000A78_00000A77_00000A76),
      .INIT_31(256'h00000773_00000772_00000771_00000770_0000076F_0000076E_0000076D_0000076C),
      .INIT_32(256'h000008B3_000008A9_00000863_00000859_00000813_00000809_000007C3_000007B9),
      .INIT_33(256'h000009F3_000009E9_000009A3_00000999_00000953_00000949_00000903_000008F9),
      .INIT_34(256'h00000A8E_00000A8D_00000A8C_00000A8B_00000A8A_00000A89_00000A43_00000A39),
      .INIT_35(256'h00000D29_00000D28_00000D27_00000A93_00000A92_00000A91_00000A90_00000A8F),
      .INIT_36(256'h00000D31_00000D30_00000D2F_00000D2E_00000D2D_00000D2C_00000D2B_00000D2A),
      .INIT_37(256'h00000E71_00000E67_00000E21_00000E17_00000DD1_00000DC7_00000D81_00000D77),
      .INIT_38(256'h00000FB1_00000FA7_00000F61_00000F57_00000F11_00000F07_00000EC1_00000EB7),
      .INIT_39(256'h0000104C_0000104B_0000104A_00001049_00001048_00001047_00001001_00000FF7),
      .INIT_3A(256'h00000D42_00000D41_00000D40_00001051_00001050_0000104F_0000104E_0000104D),
      .INIT_3B(256'h00000D4A_00000D49_00000D48_00000D47_00000D46_00000D45_00000D44_00000D43),
      .INIT_3C(256'h00000E8A_00000E80_00000E3A_00000E30_00000DEA_00000DE0_00000D9A_00000D90),
      .INIT_3D(256'h00000FCA_00000FC0_00000F7A_00000F70_00000F2A_00000F20_00000EDA_00000ED0),
      .INIT_3E(256'h00001065_00001064_00001063_00001062_00001061_00001060_0000101A_00001010),
      .INIT_3F(256'h00000D5B_00000D5A_00000D59_0000106A_00001069_00001068_00001067_00001066),


      // The next set of INITP_xx are for the parity bits
      // Address 0 to 127
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 128 to 255
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 256 to 383
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 384 to 511
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) 
 DM_inst1 (
      .DO(dm_a),      // 32-bit Data Output
      .DOP(),    // 4-bit parity Output
      .ADDR(addr_in[8:0]),  // 9-bit Address Input
      .CLK(clk),    // Clock
      .DI(fw_dm),      // 32-bit Data Input
      .DIP(4'd0),    // 4-bit parity Input
      .EN(d_enbl_a),      // RAM Enable Input
      .SSR(rst),    // Synchronous Set/Reset Input
      .WE(ctl3)       // Write Enable Input
   );

 // End of RAMB16_S36_inst instantiatio
 				
//  RAMB16_S36 : In order to incorporate this function into the design,
//   Verilog   : the following instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB16_S36_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

// RAMB16_S36: 512 x 32 + 4 Parity bits Single-Port RAM
//             Spartan-3E
// Xilinx HDL Language Template, version 12.1
RAMB16_S36 #(
      .INIT(36'h000000000),  // Value of output RAM registers at startup
      .SRVAL(36'h000000000), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 127
      // Address 0 to 127
      .INIT_00(256'h00000D63_00000D62_00000D61_00000D60_00000D5F_00000D5E_00000D5D_00000D5C),
      .INIT_01(256'h00000EA3_00000E99_00000E53_00000E49_00000E03_00000DF9_00000DB3_00000DA9),
      .INIT_02(256'h00000FE3_00000FD9_00000F93_00000F89_00000F43_00000F39_00000EF3_00000EE9),
      .INIT_03(256'h0000107E_0000107D_0000107C_0000107B_0000107A_00001079_00001033_00001029),
      .INIT_04(256'h00000000_00000000_00000000_00001083_00001082_00001081_00001080_0000107F),
      .INIT_05(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_06(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_07(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_08(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_09(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_0F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 128 to 255
      .INIT_10(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_11(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_12(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_13(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_14(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_15(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_16(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_17(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_18(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_19(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_1F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 256 to 383
      .INIT_20(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_21(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_22(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_23(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_24(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_25(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_26(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_27(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_28(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_29(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_2F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      // Address 384 to 511
      .INIT_30(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_31(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_32(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_33(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_34(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_35(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_36(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_37(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_38(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_39(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3A(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3B(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3C(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3D(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3E(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),
      .INIT_3F(256'h00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000),

      // The next set of INITP_xx are for the parity bits
      // Address 0 to 127
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 128 to 255
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 256 to 383
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 384 to 511
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) 
 DM_inst2 (
      .DO(dm_b),      // 32-bit Data Output
      .DOP(),    // 4-bit parity Output
      .ADDR(addr_in[8:0]),  // 9-bit Address Input
      .CLK(clk),    // Clock
      .DI(fw_dm),      // 32-bit Data Input
      .DIP(4'd0),    // 4-bit parity Input
      .EN(map_and),      // RAM Enable Input
      .SSR(rst),    // Synchronous Set/Reset Input
      .WE(ctl3)       // Write Enable Input
   );

 // End of RAMB16_S36_inst instantiatio
 //////////MAP Register load enable////
 assign map_e = (addr_in[9:0] == 700);
 ///////////And Gate /////////
 always@(*)
 map_and = (d_enbl_b) & ~(map_e);
  always@(posedge clk)
    begin
	 if(rst)
	    r_map <= 0;
    else if((interrupt1)|(map_e))
       r_map <= {interrupt1,23'd0,key_code1};	 
	 else
	    r_map <= r_map;
	 end
////////Mux1/////
	always@(*)
  begin
  case(d_enbl_b)
    1'd0:  dm_out1 = dm_a;
    1'd1: dm_out1 = dm_b;
    
  endcase
end
/////////Mux2////////
always@(*)
  begin
  case(map_e)
    1'd0:  dm_out = dm_out1;
    1'd1: dm_out = r_map;
    
  endcase
end		
 //dmmm endd
  //MUX for ALU
  always@(*)
  begin
  case(ctl8)
    1'd0: data2_alu_in={{15{inst_out[16]}},inst_out[16:0]};
    1'd1: data2_alu_in=reg_out2;
    
  endcase
end		

//Pipelining before ALU

//Inst register 
always@(posedge clk)
   begin
     if(rst)
      inst_r_1 <=#1 0;
     else
       inst_r_1 <=#1 inst_out;
   end  

//Reg File Data 1 Register
always@(posedge clk)
   begin
     if(rst)
      reg_d01 <=#1 0;
     else
       reg_d01 <=#1 reg_out1;
   end

//Reg File MUX of Data 2+ Inst data Register
always@(posedge clk)
   begin
     if(rst)
      mux_d02 <= #1 0;
     else
       mux_d02 <= #1 data2_alu_in;
   end

// 1st Register For CTL2
always@(posedge clk)
   begin
     if(rst)
      ctl2_1 <= #1 0;
     else
       ctl2_1 <= #1 ctl2;
   end   

// 1st Register For CTL7
always@(posedge clk)
   begin
     if(rst)
      ctl7_1 <= #1 0;
     else
      ctl7_1 <= #1 ctl7;
   end  

// 1st Register For CTL1
always@(posedge clk)
   begin
     if(rst)
      ctl1_1 <= #1 0;
     else
      ctl1_1 <= #1 ctl1;
   end 
   
// 1st Register For lui
always@(posedge clk)
   begin
     if(rst)
      lui_1 <= #1 0;
     else
      lui_1 <= #1 lui;
   end 
   
// 1st Register For lli
always@(posedge clk)
   begin
     if(rst)
      lli_1 <= #1 0;
     else
      lli_1 <= #1 lli;
   end 
  
// end of Pipelining before ALU

//Mux's for Forwarding(Read After Write )

//Mux data_1 Select Line
assign sel_md1=(inst_r_1[21:17]==inst_r_2[26:22]);
//Mux data_1 
  always@(*)
  begin
  case(sel_md1)
    1'd0: fw_d1=reg_d01;
    1'd1: fw_d1=mux_alu_o;
    
  endcase
end	

//Mux data_2 Select Line
assign sel_md2=(inst_r_1[16:12]==inst_r_2[26:22]);
//Mux data_2 
  always@(*)
  begin
  case(sel_md2)
    1'd0: fw_d2=mux_d02;
    1'd1: fw_d2=mux_alu_o;
    
  endcase
end
//end forwarding

//ALU Unit          
ALU inst3(
 .clk(clk),
 .rst(rst),
 .sel_m1(inst_r_1[28:27]),
 .data_1(fw_d1),
 .data_2(fw_d2),
 .data_out(data_alu_out)
  ); 
  
endmodule