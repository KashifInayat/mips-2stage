`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:55:43 12/27/2012 
// Design Name: 
// Module Name:    logic 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
/////////////////////////////////////////////////////////////////////////////////////////////////////////
module logic_game(
input clk,
input reset,
input [12:0] b_add,
output reg[7:0] vga_clr
    );
wire en_1;
wire en_2;
wire en_3;
wire [7:0]out_1;
wire [7:0]out_2;
wire [7:0]out_3;
//////////Enable of Block RAM 1///////////
assign en_1= (b_add[13:12]==2'b00);
//////////Enable of Block RAM 1///////////
assign en_2= (b_add[13:12]==2'b01);
//////////Enable of Block RAM 1///////////
assign en_3= (b_add[13:12]==2'b10);


//  RAMB16_S9_S9 : In order to incorporate this function into the design,
//    Verilog    : the following instance declaration needs to be placed
//   instance    : in the body of the design code.  The instance name
//  declaration  : (RAMB16_S9_S9_inst) and/or the port declarations within the
//     code      : parenthesis may be changed to properly reference and
//               : connect this function to the design.  All inputs
//               : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB16_S9_S9: 2k x 8 + 1 Parity bit Dual-Port RAM
   //               Spartan-3E
   // Xilinx HDL Language Template, version 12.1

   RAMB16_S9_S9 #(
      .INIT_A(9'h000),  // Value of output RAM registers on Port A at startup
      .INIT_B(9'h000),  // Value of output RAM registers on Port B at startup
      .SRVAL_A(9'h000), // Port A output value upon SSR assertion
      .SRVAL_B(9'h000), // Port B output value upon SSR assertion
      .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .SIM_COLLISION_CHECK("ALL"), // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 511
		                
      .INIT_00(256'hE0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),
      .INIT_01(256'hE0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),
      .INIT_02(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),
      .INIT_03(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_04(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_05(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_06(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_07(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_08(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_09(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_0A(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_0B(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_0E(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_0F(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      // Address 512 to 1023
      .INIT_10(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_11(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_12(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_13(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_14(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),//640,
      .INIT_15(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_16(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_17(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_18(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_19(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_1A(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_1D(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),//928
      .INIT_1E(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),//31
      .INIT_1F(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_992),
      // Address 1024 to 1535
      .INIT_20(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_21(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_22(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_23(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),//1120(36)
      .INIT_24(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_25(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_26(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_27(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),//(40)
      .INIT_28(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),//1280
      .INIT_29(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_2C(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_2D(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_2E(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2F(256'hE0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),//(48)(1504)
      // Address 1536 to 2047
      .INIT_30(256'hE0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),
      .INIT_31(256'h00_00_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),
      .INIT_32(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_33(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_34(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),//(53)
      .INIT_35(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_36(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_37(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_38(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_39(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_3B(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_3C(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_3D(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
		
		
		
		
      // The next set of INITP_xx are for the parity bits
      // Address 0 to 511
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 512 to 1023
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 1024 to 1535
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 1536 to 2047
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S9_S9_inst1 (
      .DOA(out_1),      // Port A 8-bit Data Output
      .DOB(DOB),      // Port B 8-bit Data Output
      .DOPA(DOPA),    // Port A 1-bit Parity Output
      .DOPB(DOPB),    // Port B 1-bit Parity Output
      .ADDRA(b_add[10:0]),  // Port A 11-bit Address Input
      .ADDRB(ADDRB),  // Port B 11-bit Address Input
      .CLKA(clk),    // Port A Clock
      .CLKB(CLKB),    // Port B Clock
      .DIA(8'd0),      // Port A 8-bit Data Input
      .DIB(DIB),      // Port B 8-bit Data Input
      .DIPA(DIPA),    // Port A 1-bit parity Input
      .DIPB(DIPB),    // Port-B 1-bit parity Input
      .ENA(en_1),      // Port A RAM Enable Input
      .ENB(ENB),      // Port B RAM Enable Input
      .SSRA(reset),    // Port A Synchronous Set/Reset Input
      .SSRB(SSRB),    // Port B Synchronous Set/Reset Input
      .WEA(1'd0),      // Port A Write Enable Input
      .WEB(WEB)       // Port B Write Enable Input
   );

   // End of RAMB16_S9_S9_inst instantiation
						
						
						
						
						
						
///////////////////////////// 2nd /////////////////////////////////////////////////////						

//  RAMB16_S9_S9 : In order to incorporate this function into the design,
//    Verilog    : the following instance declaration needs to be placed
//   instance    : in the body of the design code.  The instance name
//  declaration  : (RAMB16_S9_S9_inst) and/or the port declarations within the
//     code      : parenthesis may be changed to properly reference and
//               : connect this function to the design.  All inputs
//               : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB16_S9_S9: 2k x 8 + 1 Parity bit Dual-Port RAM
   //               Spartan-3E
   // Xilinx HDL Language Template, version 12.1

   RAMB16_S9_S9 #(
      .INIT_A(9'h000),  // Value of output RAM registers on Port A at startup
      .INIT_B(9'h000),  // Value of output RAM registers on Port B at startup
      .SRVAL_A(9'h000), // Port A output value upon SSR assertion
      .SRVAL_B(9'h000), // Port B output value upon SSR assertion
      .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .SIM_COLLISION_CHECK("ALL"), // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 511

      .INIT_00(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),//(2048)(65)
      .INIT_01(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_02(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_03(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_04(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_05(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_06(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_07(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_08(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_09(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_0A(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_0B(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_0C(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_0F(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      // Address 512 to 1023
      .INIT_10(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_11(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_12(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_13(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_14(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_15(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_16(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_17(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_18(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_19(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),//(90)
      .INIT_1A(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_1B(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_1E(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_1F(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),//(96)
      // Address 1024 to 1535
      .INIT_20(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),//(3072)
      .INIT_21(256'hE0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),//(3104)
      .INIT_22(256'hE0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),
      .INIT_23(256'h00_00_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),
      .INIT_24(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),//(3200)
      .INIT_25(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_26(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_27(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_28(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_29(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_2A(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_2D(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),//110)
      .INIT_2E(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_2F(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      // Address 1536 to 2047
      .INIT_30(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_31(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_32(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_33(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_34(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_35(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_36(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_37(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_38(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_39(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_3C(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_3D(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_3E(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),//(128)
// The next set of INITP_xx are for the parity bits
      // Address 0 to 511
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 512 to 1023
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 1024 to 1535
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 1536 to 2047
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S9_S9_inst2 (
      .DOA(out_2),      // Port A 8-bit Data Output
      .DOB(DOB),      // Port B 8-bit Data Output
      .DOPA(DOPA),    // Port A 1-bit Parity Output
      .DOPB(DOPB),    // Port B 1-bit Parity Output
      .ADDRA(b_add[10:0]),  // Port A 11-bit Address Input
      .ADDRB(ADDRB),  // Port B 11-bit Address Input
      .CLKA(clk),    // Port A Clock
      .CLKB(CLKB),    // Port B Clock
      .DIA(8'd0),      // Port A 8-bit Data Input
      .DIB(DIB),      // Port B 8-bit Data Input
      .DIPA(DIPA),    // Port A 1-bit parity Input
      .DIPB(DIPB),    // Port-B 1-bit parity Input
      .ENA(en_2),      // Port A RAM Enable Input
      .ENB(ENB),      // Port B RAM Enable Input
      .SSRA(reset),    // Port A Synchronous Set/Reset Input
      .SSRB(SSRB),    // Port B Synchronous Set/Reset Input
      .WEA(1'd0),      // Port A Write Enable Input
      .WEB(WEB)       // Port B Write Enable Input
		);

   // End of RAMB16_S9_S9_inst instantiation
	
	////////////////////////////////////////  3rd  ////////////////////////////////////////////////
	
//  RAMB16_S9_S9 : In order to incorporate this function into the design,
//    Verilog    : the following instance declaration needs to be placed
//   instance    : in the body of the design code.  The instance name
//  declaration  : (RAMB16_S9_S9_inst) and/or the port declarations within the
//     code      : parenthesis may be changed to properly reference and
//               : connect this function to the design.  All inputs
//               : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB16_S9_S9: 2k x 8 + 1 Parity bit Dual-Port RAM
   //               Spartan-3E
   // Xilinx HDL Language Template, version 12.1

   RAMB16_S9_S9 #(
      .INIT_A(9'h000),  // Value of output RAM registers on Port A at startup
      .INIT_B(9'h000),  // Value of output RAM registers on Port B at startup
      .SRVAL_A(9'h000), // Port A output value upon SSR assertion
      .SRVAL_B(9'h000), // Port B output value upon SSR assertion
      .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .SIM_COLLISION_CHECK("ALL"), // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 511
      
      .INIT_00(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_01(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_02(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_03(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_04(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_05(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_06(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_07(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_08(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_09(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      .INIT_0B(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),
      .INIT_0C(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_0D(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_0F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00),
      // Address 512 to 1023
      .INIT_10(256'h00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00),//(4608)
      .INIT_11(256'h00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_E0),
      .INIT_12(256'h00_00_00_00_00_00_00_00_00_00_00_00_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_13(256'hE0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),//(4704)
      .INIT_14(256'hE0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),
      .INIT_15(256'h00_00_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0_E0),//(150)
      .INIT_16(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_17(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_18(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_19(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_1F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      // Address 1024 to 1535
      .INIT_20(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_21(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_22(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_23(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_24(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_25(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_26(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_27(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_28(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_29(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_2F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      // Address 1536 to 2047
      .INIT_30(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_31(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_32(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_33(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_34(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_35(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_36(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_37(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_38(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_39(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3A(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3B(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3C(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3D(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3E(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),
      .INIT_3F(256'h00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00_00),

      // The next set of INITP_xx are for the parity bits
      // Address 0 to 511
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 512 to 1023
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 1024 to 1535
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 1536 to 2047
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S9_S9_inst3 (
      .DOA(out_3),      // Port A 8-bit Data Output
      .DOB(DOB),      // Port B 8-bit Data Output
      .DOPA(DOPA),    // Port A 1-bit Parity Output
      .DOPB(DOPB),    // Port B 1-bit Parity Output
      .ADDRA(b_add[10:0]),  // Port A 11-bit Address Input
      .ADDRB(ADDRB),  // Port B 11-bit Address Input
      .CLKA(clk),    // Port A Clock
      .CLKB(CLKB),    // Port B Clock
      .DIA(8'd0),      // Port A 8-bit Data Input
      .DIB(DIB),      // Port B 8-bit Data Input
      .DIPA(DIPA),    // Port A 1-bit parity Input
      .DIPB(DIPB),    // Port-B 1-bit parity Input
      .ENA(en_3),      // Port A RAM Enable Input
      .ENB(ENB),      // Port B RAM Enable Input
      .SSRA(reset),    // Port A Synchronous Set/Reset Input
      .SSRB(SSRB),    // Port B Synchronous Set/Reset Input
      .WEA(1'd0),      // Port A Write Enable Input
      .WEB(WEB)       // Port B Write Enable Input
   );

   // End of RAMB16_S9_S9_inst instantiation
always@(*)
begin
   case(b_ad[12:11])
   2'd0: vga_clr= out_1;
   2'd1: vga_clr= out_2;
   2'd2: vga_clr= out_3;
   2'd3: vga_clr= 0;
   endcase
end						